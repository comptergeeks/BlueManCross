module DE1_SoC (HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, KEY, LEDR, SW,
                CLOCK_50, VGA_R, VGA_G, VGA_B, VGA_BLANK_N, VGA_CLK, VGA_HS, VGA_SYNC_N, VGA_VS);
    output logic [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;
    output logic [9:0] LEDR;
    input logic [3:0] KEY;
    input logic [9:0] SW;
    input CLOCK_50;
    output [7:0] VGA_R;
    output [7:0] VGA_G;
    output [7:0] VGA_B;
    output VGA_BLANK_N;
    output VGA_CLK;
    output VGA_HS;
    output VGA_SYNC_N;
    output VGA_VS;
    logic [9:0] x;
    logic [8:0] y;
    logic [7:0] r, g, b;

    video_driver #(.WIDTH(640), .HEIGHT(480))
        v1 (.CLOCK_50, .reset(SW[9]), .x, .y, .r, .g, .b,
            .VGA_R, .VGA_G, .VGA_B, .VGA_BLANK_N,
            .VGA_CLK, .VGA_HS, .VGA_SYNC_N, .VGA_VS,
            .start(SW[0]), .KEY(KEY), .SW(SW)
        );

    always_ff @(posedge CLOCK_50) begin
        r <= SW[7:0];
        g <= x[7:0];
        b <= y[7:0];
    end
    
    assign HEX0 = '1;
    assign HEX1 = '1;
    assign HEX2 = '1;
    assign HEX3 = '1;
    assign HEX4 = '1;
    assign HEX5 = '1;
    
endmodule